library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;

entity fsk_timer is
    port (
        reset_n     : in    std_logic;
        clk         : in    std_logic
    );
end fsk_timer;

architecture behaviour of fsk_timer is

-- Constants

-- Signals

begin
end architecture behaviour;
